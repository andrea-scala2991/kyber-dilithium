`timescale 1ns / 1ps

module twiddle_ROM (
    input  logic        clk,
    input  logic [7:0]  addr,   // 0-255
    output logic [11:0] dout
);

    // Internal signal for combinational lookup
    logic [11:0] rom_data;

    always_comb begin
        unique case (addr)
            8'd0:   rom_data = 12'd1;
            8'd1:   rom_data = 12'd3328;
            8'd2:   rom_data = 12'd1600;
            8'd3:   rom_data = 12'd1729;
            8'd4:   rom_data = 12'd40;
            8'd5:   rom_data = 12'd3289;
            8'd6:   rom_data = 12'd749;
            8'd7:   rom_data = 12'd2580;
            8'd8:   rom_data = 12'd2481;
            8'd9:   rom_data = 12'd848;
            8'd10:  rom_data = 12'd1432;
            8'd11:  rom_data = 12'd1897;
            8'd12:  rom_data = 12'd2699;
            8'd13:  rom_data = 12'd630;
            8'd14:  rom_data = 12'd687;
            8'd15:  rom_data = 12'd2642;
            8'd16:  rom_data = 12'd1583;
            8'd17:  rom_data = 12'd1746;
            8'd18:  rom_data = 12'd2760;
            8'd19:  rom_data = 12'd569;
            8'd20:  rom_data = 12'd69;
            8'd21:  rom_data = 12'd3260;
            8'd22:  rom_data = 12'd543;
            8'd23:  rom_data = 12'd2786;
            8'd24:  rom_data = 12'd2532;
            8'd25:  rom_data = 12'd797;
            8'd26:  rom_data = 12'd3136;
            8'd27:  rom_data = 12'd193;
            8'd28:  rom_data = 12'd1410;
            8'd29:  rom_data = 12'd1919;
            8'd30:  rom_data = 12'd2267;
            8'd31:  rom_data = 12'd1062;
            8'd32:  rom_data = 12'd2508;
            8'd33:  rom_data = 12'd821;
            8'd34:  rom_data = 12'd1355;
            8'd35:  rom_data = 12'd1974;
            8'd36:  rom_data = 12'd450;
            8'd37:  rom_data = 12'd2879;
            8'd38:  rom_data = 12'd936;
            8'd39:  rom_data = 12'd2393;
            8'd40:  rom_data = 12'd447;
            8'd41:  rom_data = 12'd2882;
            8'd42:  rom_data = 12'd2794;
            8'd43:  rom_data = 12'd535;
            8'd44:  rom_data = 12'd1235;
            8'd45:  rom_data = 12'd2094;
            8'd46:  rom_data = 12'd1903;
            8'd47:  rom_data = 12'd1426;
            8'd48:  rom_data = 12'd1996;
            8'd49:  rom_data = 12'd1333;
            8'd50:  rom_data = 12'd1089;
            8'd51:  rom_data = 12'd2240;
            8'd52:  rom_data = 12'd3273;
            8'd53:  rom_data = 12'd56;
            8'd54:  rom_data = 12'd283;
            8'd55:  rom_data = 12'd3046;
            8'd56:  rom_data = 12'd1853;
            8'd57:  rom_data = 12'd1476;
            8'd58:  rom_data = 12'd1990;
            8'd59:  rom_data = 12'd1339;
            8'd60:  rom_data = 12'd882;
            8'd61:  rom_data = 12'd2447;
            8'd62:  rom_data = 12'd3033;
            8'd63:  rom_data = 12'd296;
            8'd64:  rom_data = 12'd910;
            8'd65:  rom_data = 12'd2419;
            8'd66:  rom_data = 12'd1227;
            8'd67:  rom_data = 12'd2102;
            8'd68:  rom_data = 12'd3110;
            8'd69:  rom_data = 12'd219;
            8'd70:  rom_data = 12'd2474;
            8'd71:  rom_data = 12'd855;
            8'd72:  rom_data = 12'd648;
            8'd73:  rom_data = 12'd2681;
            8'd74:  rom_data = 12'd1481;
            8'd75:  rom_data = 12'd1848;
            8'd76:  rom_data = 12'd2617;
            8'd77:  rom_data = 12'd712;
            8'd78:  rom_data = 12'd2647;
            8'd79:  rom_data = 12'd682;
            8'd80:  rom_data = 12'd2402;
            8'd81:  rom_data = 12'd927;
            8'd82:  rom_data = 12'd1534;
            8'd83:  rom_data = 12'd1795;
            8'd84:  rom_data = 12'd2868;
            8'd85:  rom_data = 12'd461;
            8'd86:  rom_data = 12'd1438;
            8'd87:  rom_data = 12'd1891;
            8'd88:  rom_data = 12'd452;
            8'd89:  rom_data = 12'd2877;
            8'd90:  rom_data = 12'd807;
            8'd91:  rom_data = 12'd2522;
            8'd92:  rom_data = 12'd1435;
            8'd93:  rom_data = 12'd1894;
            8'd94:  rom_data = 12'd2319;
            8'd95:  rom_data = 12'd1010;
            8'd96:  rom_data = 12'd1915;
            8'd97:  rom_data = 12'd1414;
            8'd98:  rom_data = 12'd1320;
            8'd99:  rom_data = 12'd2009;
            8'd100: rom_data = 12'd33;
            8'd101: rom_data = 12'd3296;
            8'd102: rom_data = 12'd2865;
            8'd103: rom_data = 12'd464;
            8'd104: rom_data = 12'd632;
            8'd105: rom_data = 12'd2697;
            8'd106: rom_data = 12'd2513;
            8'd107: rom_data = 12'd816;
            8'd108: rom_data = 12'd1977;
            8'd109: rom_data = 12'd1352;
            8'd110: rom_data = 12'd650;
            8'd111: rom_data = 12'd2679;
            8'd112: rom_data = 12'd2055;
            8'd113: rom_data = 12'd1274;
            8'd114: rom_data = 12'd2277;
            8'd115: rom_data = 12'd1052;
            8'd116: rom_data = 12'd2304;
            8'd117: rom_data = 12'd1025;
            8'd118: rom_data = 12'd1197;
            8'd119: rom_data = 12'd2132;
            8'd120: rom_data = 12'd1756;
            8'd121: rom_data = 12'd1573;
            8'd122: rom_data = 12'd3253;
            8'd123: rom_data = 12'd76;
            8'd124: rom_data = 12'd331;
            8'd125: rom_data = 12'd2998;
            8'd126: rom_data = 12'd289;
            8'd127: rom_data = 12'd3040;
            8'd128: rom_data = 12'd1;
            8'd129: rom_data = 12'd3328;
            8'd130: rom_data = 12'd1729;
            8'd131: rom_data = 12'd1600;
            8'd132: rom_data = 12'd2580;
            8'd133: rom_data = 12'd749;
            8'd134: rom_data = 12'd3289;
            8'd135: rom_data = 12'd40;
            8'd136: rom_data = 12'd2642;
            8'd137: rom_data = 12'd687;
            8'd138: rom_data = 12'd630;
            8'd139: rom_data = 12'd2699;
            8'd140: rom_data = 12'd1897;
            8'd141: rom_data = 12'd1432;
            8'd142: rom_data = 12'd848;
            8'd143: rom_data = 12'd2481;
            8'd144: rom_data = 12'd1062;
            8'd145: rom_data = 12'd2267;
            8'd146: rom_data = 12'd1919;
            8'd147: rom_data = 12'd1410;
            8'd148: rom_data = 12'd193;
            8'd149: rom_data = 12'd3136;
            8'd150: rom_data = 12'd797;
            8'd151: rom_data = 12'd2532;
            8'd152: rom_data = 12'd2786;
            8'd153: rom_data = 12'd543;
            8'd154: rom_data = 12'd3260;
            8'd155: rom_data = 12'd69;
            8'd156: rom_data = 12'd569;
            8'd157: rom_data = 12'd2760;
            8'd158: rom_data = 12'd1746;
            8'd159: rom_data = 12'd1583;
            8'd160: rom_data = 12'd296;
            8'd161: rom_data = 12'd3033;
            8'd162: rom_data = 12'd2447;
            8'd163: rom_data = 12'd882;
            8'd164: rom_data = 12'd1339;
            8'd165: rom_data = 12'd1990;
            8'd166: rom_data = 12'd1476;
            8'd167: rom_data = 12'd1853;
            8'd168: rom_data = 12'd3046;
            8'd169: rom_data = 12'd283;
            8'd170: rom_data = 12'd56;
            8'd171: rom_data = 12'd3273;
            8'd172: rom_data = 12'd2240;
            8'd173: rom_data = 12'd1089;
            8'd174: rom_data = 12'd1333;
            8'd175: rom_data = 12'd1996;
            8'd176: rom_data = 12'd1426;
            8'd177: rom_data = 12'd1903;
            8'd178: rom_data = 12'd2094;
            8'd179: rom_data = 12'd1235;
            8'd180: rom_data = 12'd535;
            8'd181: rom_data = 12'd2794;
            8'd182: rom_data = 12'd2882;
            8'd183: rom_data = 12'd447;
            8'd184: rom_data = 12'd2393;
            8'd185: rom_data = 12'd936;
            8'd186: rom_data = 12'd2879;
            8'd187: rom_data = 12'd450;
            8'd188: rom_data = 12'd1974;
            8'd189: rom_data = 12'd1355;
            8'd190: rom_data = 12'd821;
            8'd191: rom_data = 12'd2508;
            8'd192: rom_data = 12'd3040;
            8'd193: rom_data = 12'd289;
            8'd194: rom_data = 12'd2998;
            8'd195: rom_data = 12'd331;
            8'd196: rom_data = 12'd76;
            8'd197: rom_data = 12'd3253;
            8'd198: rom_data = 12'd1573;
            8'd199: rom_data = 12'd1756;
            8'd200: rom_data = 12'd2132;
            8'd201: rom_data = 12'd1197;
            8'd202: rom_data = 12'd1025;
            8'd203: rom_data = 12'd2304;
            8'd204: rom_data = 12'd1052;
            8'd205: rom_data = 12'd2277;
            8'd206: rom_data = 12'd1274;
            8'd207: rom_data = 12'd2055;
            8'd208: rom_data = 12'd2679;
            8'd209: rom_data = 12'd650;
            8'd210: rom_data = 12'd1352;
            8'd211: rom_data = 12'd1977;
            8'd212: rom_data = 12'd816;
            8'd213: rom_data = 12'd2513;
            8'd214: rom_data = 12'd2697;
            8'd215: rom_data = 12'd632;
            8'd216: rom_data = 12'd464;
            8'd217: rom_data = 12'd2865;
            8'd218: rom_data = 12'd3296;
            8'd219: rom_data = 12'd33;
            8'd220: rom_data = 12'd2009;
            8'd221: rom_data = 12'd1320;
            8'd222: rom_data = 12'd1414;
            8'd223: rom_data = 12'd1915;
            8'd224: rom_data = 12'd1010;
            8'd225: rom_data = 12'd2319;
            8'd226: rom_data = 12'd1894;
            8'd227: rom_data = 12'd1435;
            8'd228: rom_data = 12'd2522;
            8'd229: rom_data = 12'd807;
            8'd230: rom_data = 12'd2877;
            8'd231: rom_data = 12'd452;
            8'd232: rom_data = 12'd1891;
            8'd233: rom_data = 12'd1438;
            8'd234: rom_data = 12'd461;
            8'd235: rom_data = 12'd2868;
            8'd236: rom_data = 12'd1795;
            8'd237: rom_data = 12'd1534;
            8'd238: rom_data = 12'd927;
            8'd239: rom_data = 12'd2402;
            8'd240: rom_data = 12'd682;
            8'd241: rom_data = 12'd2647;
            8'd242: rom_data = 12'd712;
            8'd243: rom_data = 12'd2617;
            8'd244: rom_data = 12'd1848;
            8'd245: rom_data = 12'd1481;
            8'd246: rom_data = 12'd2681;
            8'd247: rom_data = 12'd648;
            8'd248: rom_data = 12'd855;
            8'd249: rom_data = 12'd2474;
            8'd250: rom_data = 12'd219;
            8'd251: rom_data = 12'd3110;
            8'd252: rom_data = 12'd2102;
            8'd253: rom_data = 12'd1227;
            8'd254: rom_data = 12'd2419;
            8'd255: rom_data = 12'd910;
            default: rom_data = 12'd0;
        endcase
    end

    // Register output (synchronous ROM)
    always_ff @(posedge clk) begin
        dout <= rom_data;
    end

endmodule
